----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:29:40 09/10/2024 
-- Design Name: 
-- Module Name:    AND_2_Vectors_4_Bits - AND_2_Vectors_4_Bits 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity NAND_2_Vectors_4_Bits is
        Port ( A : in  STD_LOGIC_VECTOR (3 downto 0);
               B : in  STD_LOGIC_VECTOR (3 downto 0);
               C : out  STD_LOGIC_VECTOR (3 downto 0));
    end NAND_2_Vectors_4_Bits;
    
architecture Behavioral of NAND_2_Vectors_4_Bits is
    begin
        C <= NOT (A and B);
end Behavioral;
